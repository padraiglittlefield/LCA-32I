module load_store_unit (
    input clk, 
    input rst
);

//TODO: Go back and make sure everything works with all types of mem instructions

load_data_queue ldq (

);

store_data_queue sdq (
    
);

endmodule
