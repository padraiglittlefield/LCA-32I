module tb_miss_status_history_register;

endmodule