module load_store_unit (
    input clk_i, 
    input rst_i,
    input flush_i,

    dispatch_lsu_if.lsu disp_if,
    execute_lsu_if.lsu exec_if,
    lsu_reorder_buffer.lsu rob_if,
    
    output mem_req_vld_o,
    output mem_req_addr_o,
    input mem_resp_vld_i,
    input mem_resp_data_i
);

//TODO: Go back and make sure everything works with all types of mem instructions
//TODO: Make sure speculative state is flushed but that unspectulative state remains. Espically with the SDQ. I think LDQ can just be lfushed
//      ^ this is mostly implemented by it needs to be double checked

    load_data_queue u_ldq (
        .clk_i(clk_i),
        .rst_i(rst_i),
        .flush_i(flush_i),
        .disp_vld_i(),
        .disp_dsq_marker_i(),
        .ldq_disp_idx_o(),
        .ldq_full_o(),
        .exec_vld_i(),
        .exec_ldq_idx_i(),
        .exec_addr_i(),
        .issue_en_i(),
        .issue_entry_o(),
        .issue_vld_o()
    );

    store_data_queue u_sdq (
        .clk_i(clk_i),
        .rst_i(rst_i),
        .flush_i(flush_i),
        .disp_vld_i(),
        .store_data_i(),
        .cmit_vld_i(),
        .cmit_idx_i(),
        .exec_vld_i(),
        .exec_addr_i(),
        .sdq_alloc_idx_o(),
        .sdq_full_o(),
        .issue_en_i(),
        .issue_entry_o(),
        .isse_vld_o(),
        .ld_vld_i(),
        .ld_addr_i(),
        .ld_sdq_marker_i(),
        .ld_hit_o(),
        .ld_data_o()
    );

   cache_controller u_cache_controller (
    .clk_i(clk_i),
    .rst_i(rst_i),
    .flush_i(flush_i),
    .lsu_req_vld_i(),
    .lsu_req_wr_rd_i(),
    .lsu_req_addr_i(),
    .lsu_req_data_i(),
    .lsu_req_rob_idx_i(), 
    .mem_req_vld_o(),
    .mem_req_addr_o(),
    .mem_resp_vld_i(),
    .mem_resp_data_i(), 
    .mem_wb_vld_o(),
    .mem_wb_data_o(),
    .cmt_ld_vld_o(),
    .cmt_ld_data_o(),
    .cmt_rob_idx_o(),
    .stall_controller_o()
);  


// main_memory_interface u_mmu ( // Going to move this to Chip Top instead of inside the PIPELINE

// );

endmodule
