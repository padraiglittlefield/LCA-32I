`timescale 1ns/1ns

import CORE_PKG::*;

module register_read (
    input clk,
    input rst,
    scheduler_reg_read_if sched_if,
    
);
    


endmodule