module agu();
endmodule