module load_store_unit (
    input clk, 
    input rst
);



load_data_queue ldq (

);

store_data_queue sdq (
    
);

endmodule
