module store_data_queue(
    input clk,
    input rst
);

endmodule