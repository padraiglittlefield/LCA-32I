module load_store_unit (
    input clk, 
    input rst
);

//TODO: Go back and make sure everything works with all types of mem instructions

load_data_queue u_ldq (

);

store_data_queue u_sdq (
    
);

cache_controller u_cache_controller(

);



// main_memory_interface u_mmu (

// );

endmodule
