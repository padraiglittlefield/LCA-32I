`timescale 1ns/1ns


module fwrd_unit (
    
);

endmodule
